`timescale 1ns/1ns
module TotalALU( clk, dataA, dataB, Signal, control, Output, reset );
input reset ;
input clk ;
input[2:0] control ;
input [31:0] dataA ;
input [31:0] dataB ;
input [5:0] Signal ;
output [31:0] Output ;

//   Signal ( 6-bits)?
//   AND  : 36
//   OR   : 37
//   ADD  : 32
//   SUB  : 34
//   SLL  : 0
//   SLT  : 42
//   MULTU : 25

wire [31:0] temp ;
wire Cout ;
parameter AND = 6'b100100;
parameter OR  = 6'b100101;
parameter ADD = 6'b100000;
parameter SUB = 6'b100010;
parameter SLT = 6'b101010;

parameter SLL = 6'b000000;

parameter MULTU= 6'b011001;
parameter MFHI= 6'b010000;
parameter MFLO= 6'b010010;
/*
�w�q�U�ذT��
*/
//============================
wire [5:0]  SignaltoALU ;
wire [5:0]  SignaltoSHT ;
wire [5:0]  SignaltoMUL ;
wire [5:0]  SignaltoMUX ;
wire [31:0] ALUOut, HiOut, LoOut, ShifterOut ;
wire [31:0] dataOut ;
wire [63:0] MulAns ;
/*
�w�q�U�ر��u
*/
//============================


ALUControl ALUControl( .clk(clk), .Signal(Signal), .SignaltoALU(SignaltoALU), .SignaltoSHT(SignaltoSHT), .SignaltoMUL(SignaltoMUL), .SignaltoMUX(SignaltoMUX) );
ALU alu( .dataA(dataA), .dataB(dataB), .control(control), .sum(ALUOut), .Cout(Cout) );
multiplier multiplier( .multiplicand(dataA), .multiplier(dataB), .clk(clk), .dataout(MulAns), .reset(reset) ) ;
shifter shifter( .datain(dataA), .shiftnum(dataB), .dataout(ShifterOut) ) ;
HiLo HiLo( .clk(clk), .MulAns(MulAns), .HiOut(HiOut), .LoOut(LoOut), .reset(reset) );
MUX MUX( .ALUOut(ALUOut), .HiOut(HiOut), .LoOut(LoOut), .Shifter(ShifterOut), .Cout(Cout), .Signal(SignaltoMUX), .dataOut(dataOut) );


/*
�إߦU��module
*/
assign Output = dataOut ;


endmodule